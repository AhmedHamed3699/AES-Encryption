module InverseSbox(sbox_byte,byte);
input  [7:0] sbox_byte; 
output reg [7:0] byte;

 always@(*)
 begin  
    case(sbox_byte)
				8'h00:byte =8'h52;
				8'h01:byte =8'h09;
				8'h02:byte =8'h6a;
				8'h03:byte =8'hd5;
				8'h04:byte =8'h30;
				8'h05:byte =8'h36;
				8'h06:byte =8'ha5;
				8'h07:byte =8'h38;
				8'h08:byte =8'hbf;
				8'h09:byte =8'h40;
				8'h0a:byte =8'ha3;
				8'h0b:byte =8'h9e;
				8'h0c:byte =8'h81;
				8'h0d:byte =8'hf3;
				8'h0e:byte =8'hd7;
				8'h0f:byte =8'hfb;
				8'h10:byte =8'h7c;
				8'h11:byte =8'he3;
				8'h12:byte =8'h39;
				8'h13:byte =8'h82;
				8'h14:byte =8'h9b;
				8'h15:byte =8'h2f;
				8'h16:byte =8'hff;
				8'h17:byte =8'h87;
				8'h18:byte =8'h34;
				8'h19:byte =8'h8e;
				8'h1a:byte =8'h43;
				8'h1b:byte =8'h44;
				8'h1c:byte =8'hc4;
				8'h1d:byte =8'hde;
				8'h1e:byte =8'he9;
				8'h1f:byte =8'hcb;
				8'h20:byte =8'h54;
				8'h21:byte =8'h7b;
				8'h22:byte =8'h94;
				8'h23:byte =8'h32;
				8'h24:byte =8'ha6;
				8'h25:byte =8'hc2;
				8'h26:byte =8'h23;
				8'h27:byte =8'h3d;
				8'h28:byte =8'hee;
				8'h29:byte =8'h4c;
				8'h2a:byte =8'h95;
				8'h2b:byte =8'h0b;
				8'h2c:byte =8'h42;
				8'h2d:byte =8'hfa;
				8'h2e:byte =8'hc3;
				8'h2f:byte =8'h4e;
				8'h30:byte =8'h08;
				8'h31:byte =8'h2e;
				8'h32:byte =8'ha1;
				8'h33:byte =8'h66;
				8'h34:byte =8'h28;
				8'h35:byte =8'hd9;
				8'h36:byte =8'h24;
				8'h37:byte =8'hb2;
				8'h38:byte =8'h76;
				8'h39:byte =8'h5b;
				8'h3a:byte =8'ha2;
				8'h3b:byte =8'h49;
				8'h3c:byte =8'h6d;
				8'h3d:byte =8'h8b;
				8'h3e:byte =8'hd1;
				8'h3f:byte =8'h25;
				8'h40:byte =8'h72;
				8'h41:byte =8'hf8;
				8'h42:byte =8'hf6;
				8'h43:byte =8'h64;
				8'h44:byte =8'h86;
				8'h45:byte =8'h68;
				8'h46:byte =8'h98;
				8'h47:byte =8'h16;
				8'h48:byte =8'hd4;
				8'h49:byte =8'ha4;
				8'h4a:byte =8'h5c;
				8'h4b:byte =8'hcc;
				8'h4c:byte =8'h5d;
				8'h4d:byte =8'h65;
				8'h4e:byte =8'hb6;
				8'h4f:byte =8'h92;
				8'h50:byte =8'h6c;
				8'h51:byte =8'h70;
				8'h52:byte =8'h48;
				8'h53:byte =8'h50;
				8'h54:byte =8'hfd;
				8'h55:byte =8'hed;
				8'h56:byte =8'hb9;
				8'h57:byte =8'hda;
				8'h58:byte =8'h5e;
				8'h59:byte =8'h15;
				8'h5a:byte =8'h46;
				8'h5b:byte =8'h57;
				8'h5c:byte =8'ha7;
				8'h5d:byte =8'h8d;
				8'h5e:byte =8'h9d;
				8'h5f:byte =8'h84;
				8'h60:byte =8'h90;
				8'h61:byte =8'hd8;
				8'h62:byte =8'hab;
				8'h63:byte =8'h00;
				8'h64:byte =8'h8c;
				8'h65:byte =8'hbc;
				8'h66:byte =8'hd3;
				8'h67:byte =8'h0a;
				8'h68:byte =8'hf7;
				8'h69:byte =8'he4;
				8'h6a:byte =8'h58;
				8'h6b:byte =8'h05;
				8'h6c:byte =8'hb8;
				8'h6d:byte =8'hb3;
				8'h6e:byte =8'h45;
				8'h6f:byte =8'h06;
				8'h70:byte =8'hd0;
				8'h71:byte =8'h2c;
				8'h72:byte =8'h1e;
				8'h73:byte =8'h8f;
				8'h74:byte =8'hca;
				8'h75:byte =8'h3f;
				8'h76:byte =8'h0f;
				8'h77:byte =8'h02;
				8'h78:byte =8'hc1;
				8'h79:byte =8'haf;
				8'h7a:byte =8'hbd;
				8'h7b:byte =8'h03;
				8'h7c:byte =8'h01;
				8'h7d:byte =8'h13;
				8'h7e:byte =8'h8a;
				8'h7f:byte =8'h6b;
				8'h80:byte =8'h3a;
				8'h81:byte =8'h91;
				8'h82:byte =8'h11;
				8'h83:byte =8'h41;
				8'h84:byte =8'h4f;
				8'h85:byte =8'h67;
				8'h86:byte =8'hdc;
				8'h87:byte =8'hea;
				8'h88:byte =8'h97;
				8'h89:byte =8'hf2;
				8'h8a:byte =8'hcf;
				8'h8b:byte =8'hce;
				8'h8c:byte =8'hf0;
				8'h8d:byte =8'hb4;
				8'h8e:byte =8'he6;
				8'h8f:byte =8'h73;
				8'h90:byte =8'h96;
				8'h91:byte =8'hac;
				8'h92:byte =8'h74;
				8'h93:byte =8'h22;
				8'h94:byte =8'he7;
				8'h95:byte =8'had;
				8'h96:byte =8'h35;
				8'h97:byte =8'h85;
				8'h98:byte =8'he2;
				8'h99:byte =8'hf9;
				8'h9a:byte =8'h37;
				8'h9b:byte =8'he8;
				8'h9c:byte =8'h1c;
				8'h9d:byte =8'h75;
				8'h9e:byte =8'hdf;
				8'h9f:byte =8'h6e;
				8'ha0:byte =8'h47;
				8'ha1:byte =8'hf1;
				8'ha2:byte =8'h1a;
				8'ha3:byte =8'h71;
				8'ha4:byte =8'h1d;
				8'ha5:byte =8'h29;
				8'ha6:byte =8'hc5;
				8'ha7:byte =8'h89;
				8'ha8:byte =8'h6f;
				8'ha9:byte =8'hb7;
				8'haa:byte =8'h62;
				8'hab:byte =8'h0e;
				8'hac:byte =8'haa;
				8'had:byte =8'h18;
				8'hae:byte =8'hbe;
				8'haf:byte =8'h1b;
				8'hb0:byte =8'hfc;
				8'hb1:byte =8'h56;
				8'hb2:byte =8'h3e;
				8'hb3:byte =8'h4b;
				8'hb4:byte =8'hc6;
				8'hb5:byte =8'hd2;
				8'hb6:byte =8'h79;
				8'hb7:byte =8'h20;
				8'hb8:byte =8'h9a;
				8'hb9:byte =8'hdb;
				8'hba:byte =8'hc0;
				8'hbb:byte =8'hfe;
				8'hbc:byte =8'h78;
				8'hbd:byte =8'hcd;
				8'hbe:byte =8'h5a;
				8'hbf:byte =8'hf4;
				8'hc0:byte =8'h1f;
				8'hc1:byte =8'hdd;
				8'hc2:byte =8'ha8;
				8'hc3:byte =8'h33;
				8'hc4:byte =8'h88;
				8'hc5:byte =8'h07;
				8'hc6:byte =8'hc7;
				8'hc7:byte =8'h31;
				8'hc8:byte =8'hb1;
				8'hc9:byte =8'h12;
				8'hca:byte =8'h10;
				8'hcb:byte =8'h59;
				8'hcc:byte =8'h27;
				8'hcd:byte =8'h80;
				8'hce:byte =8'hec;
				8'hcf:byte =8'h5f;
				8'hd0:byte =8'h60;
				8'hd1:byte =8'h51;
				8'hd2:byte =8'h7f;
				8'hd3:byte =8'ha9;
				8'hd4:byte =8'h19;
				8'hd5:byte =8'hb5;
				8'hd6:byte =8'h4a;
				8'hd7:byte =8'h0d;
				8'hd8:byte =8'h2d;
				8'hd9:byte =8'he5;
				8'hda:byte =8'h7a;
				8'hdb:byte =8'h9f;
				8'hdc:byte =8'h93;
				8'hdd:byte =8'hc9;
				8'hde:byte =8'h9c;
				8'hdf:byte =8'hef;
				8'he0:byte =8'ha0;
				8'he1:byte =8'he0;
				8'he2:byte =8'h3b;
				8'he3:byte =8'h4d;
				8'he4:byte =8'hae;
				8'he5:byte =8'h2a;
				8'he6:byte =8'hf5;
				8'he7:byte =8'hb0;
				8'he8:byte =8'hc8;
				8'he9:byte =8'heb;
				8'hea:byte =8'hbb;
				8'heb:byte =8'h3c;
				8'hec:byte =8'h83;
				8'hed:byte =8'h53;
				8'hee:byte =8'h99;
				8'hef:byte =8'h61;
				8'hf0:byte =8'h17;
				8'hf1:byte =8'h2b;
				8'hf2:byte =8'h04;
				8'hf3:byte =8'h7e;
				8'hf4:byte =8'hba;
				8'hf5:byte =8'h77;
				8'hf6:byte =8'hd6;
				8'hf7:byte =8'h26;
				8'hf8:byte =8'he1;
				8'hf9:byte =8'h69;
				8'hfa:byte =8'h14;
				8'hfb:byte =8'h63;
				8'hfc:byte =8'h55;
				8'hfd:byte =8'h21;
				8'hfe:byte =8'h0c;
				8'hff:byte =8'h7d;
				endcase
end

endmodule